`define zero_word 32'b0

module DataMem(
	input clk,
	input rst_n,
	
	input MemWrite,
	input MemRead,
	
	input [7:0]Address,

	input [31:0] WriteData,
	output [31:0] ReadData,
	output [31:0] IO_out
    );
	
	
	reg [31:0]ram[255:0];
	
	assign ReadData = ram[Address];
	assign IO_out = ram[0];

	always@(posedge clk)
	begin
		if(!rst_n)// for循环不知道为什么会报错，仿真暂且这样初始化
			begin
				ram[0]<=`zero_word;
				ram[1]<=`zero_word;
				ram[2]<=`zero_word;
				ram[3]<=`zero_word;
				ram[4]<=`zero_word;
				ram[5]<=`zero_word;
				ram[6]<=`zero_word;
				ram[7]<=`zero_word;
				ram[8]<=`zero_word;
				ram[9]<=`zero_word;
				ram[10]<=`zero_word;
				ram[11]<=`zero_word;
				ram[12]<=`zero_word;
				ram[13]<=`zero_word;
				ram[14]<=`zero_word;
				ram[15]<=`zero_word;
				ram[16]<=`zero_word;
				ram[17]<=`zero_word;
				ram[18]<=`zero_word;
				ram[19]<=`zero_word;
				ram[20]<=`zero_word;
				ram[21]<=`zero_word;
				ram[22]<=`zero_word;
				ram[23]<=`zero_word;
				ram[24]<=`zero_word;
				ram[25]<=`zero_word;
				ram[26]<=`zero_word;
				ram[27]<=`zero_word;
				ram[28]<=`zero_word;
				ram[29]<=`zero_word;
				ram[30]<=`zero_word;
				ram[31]<=`zero_word;
				ram[32]<=`zero_word;
				ram[33]<=`zero_word;
				ram[34]<=`zero_word;
				ram[35]<=`zero_word;
				ram[36]<=`zero_word;
				ram[37]<=`zero_word;
				ram[38]<=`zero_word;
				ram[39]<=`zero_word;
				ram[40]<=`zero_word;
				ram[41]<=`zero_word;
				ram[42]<=`zero_word;
				ram[43]<=`zero_word;
				ram[44]<=`zero_word;
				ram[45]<=`zero_word;
				ram[46]<=`zero_word;
				ram[47]<=`zero_word;
				ram[48]<=`zero_word;
				ram[49]<=`zero_word;
				ram[50]<=`zero_word;
				ram[51]<=`zero_word;
				ram[52]<=`zero_word;
				ram[53]<=`zero_word;
				ram[54]<=`zero_word;
				ram[55]<=`zero_word;
				ram[56]<=`zero_word;
				ram[57]<=`zero_word;
				ram[58]<=`zero_word;
				ram[59]<=`zero_word;
				ram[60]<=`zero_word;
				ram[61]<=`zero_word;
				ram[62]<=`zero_word;
				ram[63]<=`zero_word;
				ram[64]<=`zero_word;
				ram[65]<=`zero_word;
				ram[66]<=`zero_word;
				ram[67]<=`zero_word;
				ram[68]<=`zero_word;
				ram[69]<=`zero_word;
				ram[70]<=`zero_word;
				ram[71]<=`zero_word;
				ram[72]<=`zero_word;
				ram[73]<=`zero_word;
				ram[74]<=`zero_word;
				ram[75]<=`zero_word;
				ram[76]<=`zero_word;
				ram[77]<=`zero_word;
				ram[78]<=`zero_word;
				ram[79]<=`zero_word;
				ram[80]<=`zero_word;
				ram[81]<=`zero_word;
				ram[82]<=`zero_word;
				ram[83]<=`zero_word;
				ram[84]<=`zero_word;
				ram[85]<=`zero_word;
				ram[86]<=`zero_word;
				ram[87]<=`zero_word;
				ram[88]<=`zero_word;
				ram[89]<=`zero_word;
				ram[90]<=`zero_word;
				ram[91]<=`zero_word;
				ram[92]<=`zero_word;
				ram[93]<=`zero_word;
				ram[94]<=`zero_word;
				ram[95]<=`zero_word;
				ram[96]<=`zero_word;
				ram[97]<=`zero_word;
				ram[98]<=`zero_word;
				ram[99]<=`zero_word;
				ram[100]<=`zero_word;
				ram[101]<=`zero_word;
				ram[102]<=`zero_word;
				ram[103]<=`zero_word;
				ram[104]<=`zero_word;
				ram[105]<=`zero_word;
				ram[106]<=`zero_word;
				ram[107]<=`zero_word;
				ram[108]<=`zero_word;
				ram[109]<=`zero_word;
				ram[110]<=`zero_word;
				ram[111]<=`zero_word;
				ram[112]<=`zero_word;
				ram[113]<=`zero_word;
				ram[114]<=`zero_word;
				ram[115]<=`zero_word;
				ram[116]<=`zero_word;
				ram[117]<=`zero_word;
				ram[118]<=`zero_word;
				ram[119]<=`zero_word;
				ram[120]<=`zero_word;
				ram[121]<=`zero_word;
				ram[122]<=`zero_word;
				ram[123]<=`zero_word;
				ram[124]<=`zero_word;
				ram[125]<=`zero_word;
				ram[126]<=`zero_word;
				ram[127]<=`zero_word;
				ram[128]<=`zero_word;
				ram[129]<=`zero_word;
				ram[130]<=`zero_word;
				ram[131]<=`zero_word;
				ram[132]<=`zero_word;
				ram[133]<=`zero_word;
				ram[134]<=`zero_word;
				ram[135]<=`zero_word;
				ram[136]<=`zero_word;
				ram[137]<=`zero_word;
				ram[138]<=`zero_word;
				ram[139]<=`zero_word;
				ram[140]<=`zero_word;
				ram[141]<=`zero_word;
				ram[142]<=`zero_word;
				ram[143]<=`zero_word;
				ram[144]<=`zero_word;
				ram[145]<=`zero_word;
				ram[146]<=`zero_word;
				ram[147]<=`zero_word;
				ram[148]<=`zero_word;
				ram[149]<=`zero_word;
				ram[150]<=`zero_word;
				ram[151]<=`zero_word;
				ram[152]<=`zero_word;
				ram[153]<=`zero_word;
				ram[154]<=`zero_word;
				ram[155]<=`zero_word;
				ram[156]<=`zero_word;
				ram[157]<=`zero_word;
				ram[158]<=`zero_word;
				ram[159]<=`zero_word;
				ram[160]<=`zero_word;
				ram[161]<=`zero_word;
				ram[162]<=`zero_word;
				ram[163]<=`zero_word;
				ram[164]<=`zero_word;
				ram[165]<=`zero_word;
				ram[166]<=`zero_word;
				ram[167]<=`zero_word;
				ram[168]<=`zero_word;
				ram[169]<=`zero_word;
				ram[170]<=`zero_word;
				ram[171]<=`zero_word;
				ram[172]<=`zero_word;
				ram[173]<=`zero_word;
				ram[174]<=`zero_word;
				ram[175]<=`zero_word;
				ram[176]<=`zero_word;
				ram[177]<=`zero_word;
				ram[178]<=`zero_word;
				ram[179]<=`zero_word;
				ram[180]<=`zero_word;
				ram[181]<=`zero_word;
				ram[182]<=`zero_word;
				ram[183]<=`zero_word;
				ram[184]<=`zero_word;
				ram[185]<=`zero_word;
				ram[186]<=`zero_word;
				ram[187]<=`zero_word;
				ram[188]<=`zero_word;
				ram[189]<=`zero_word;
				ram[190]<=`zero_word;
				ram[191]<=`zero_word;
				ram[192]<=`zero_word;
				ram[193]<=`zero_word;
				ram[194]<=`zero_word;
				ram[195]<=`zero_word;
				ram[196]<=`zero_word;
				ram[197]<=`zero_word;
				ram[198]<=`zero_word;
				ram[199]<=`zero_word;
				ram[200]<=`zero_word;
				ram[201]<=`zero_word;
				ram[202]<=`zero_word;
				ram[203]<=`zero_word;
				ram[204]<=`zero_word;
				ram[205]<=`zero_word;
				ram[206]<=`zero_word;
				ram[207]<=`zero_word;
				ram[208]<=`zero_word;
				ram[209]<=`zero_word;
				ram[210]<=`zero_word;
				ram[211]<=`zero_word;
				ram[212]<=`zero_word;
				ram[213]<=`zero_word;
				ram[214]<=`zero_word;
				ram[215]<=`zero_word;
				ram[216]<=`zero_word;
				ram[217]<=`zero_word;
				ram[218]<=`zero_word;
				ram[219]<=`zero_word;
				ram[220]<=`zero_word;
				ram[221]<=`zero_word;
				ram[222]<=`zero_word;
				ram[223]<=`zero_word;
				ram[224]<=`zero_word;
				ram[225]<=`zero_word;
				ram[226]<=`zero_word;
				ram[227]<=`zero_word;
				ram[228]<=`zero_word;
				ram[229]<=`zero_word;
				ram[230]<=`zero_word;
				ram[231]<=`zero_word;
				ram[232]<=`zero_word;
				ram[233]<=`zero_word;
				ram[234]<=`zero_word;
				ram[235]<=`zero_word;
				ram[236]<=`zero_word;
				ram[237]<=`zero_word;
				ram[238]<=`zero_word;
				ram[239]<=`zero_word;
				ram[240]<=`zero_word;
				ram[241]<=`zero_word;
				ram[242]<=`zero_word;
				ram[243]<=`zero_word;
				ram[244]<=`zero_word;
				ram[245]<=`zero_word;
				ram[246]<=`zero_word;
				ram[247]<=`zero_word;
				ram[248]<=`zero_word;
				ram[249]<=`zero_word;
				ram[250]<=`zero_word;
				ram[251]<=`zero_word;
				ram[252]<=`zero_word;
				ram[253]<=`zero_word;
				ram[254]<=`zero_word;
				ram[255]<=`zero_word;
			end
		else if(MemWrite)
			ram[Address]<=WriteData;	
	end

endmodule